`define ADD  3'b000
`define ADDI 3'b001
`define MUL  3'b011
`define MULI 3'b100
`define WAIT 3'b101
`define LDSW 3'b110


