`define MOV  3'b000
`define MAC  3'b001
`define WAIT 3'b010
`define SETB 3'b011
`define SETD 3'b100
`define SETE 3'b101

