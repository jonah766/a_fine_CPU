`define MOV  3'b000
`define MAC  3'b001
`define SETB 3'b011
`define SETD 3'b100
`define SETE 3'b101
`define LDSW 3'b110
`define WAIT 3'b111


