//-----------------------------------------------------
// File Name : opcodes.sv
// Function : pMIPS instr opcode definitions
// Author: jf
//-----------------------------------------------------
//
`define NOP 6'b000000
`define ADD 6'b001010
`define SUB 6'b010011
`define ADDI 6'b011010
`define SUBI 6'b100011
`define BEQ 6'b101011
`define BNE 6'b110011
`define BGE 6'b111011
