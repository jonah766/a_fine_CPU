//-----------------------------------------------------
// File Name : opcodes.sv
// Function : pMIPS instr opcode definitions
// Author: jf
//-----------------------------------------------------
//
`define NOP  6'b000000
`define ADD  6'b000001
`define SUB  6'b000010
`define ADDI 6'b000011
`define SUBI 6'b000100
`define BEQ  6'b000101
`define BNE  6'b000110
`define BGE  6'b000111
`define BLO  6'b001000
